library work;
use work.all;
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TrafficLightContainer is
	port (clk, rst: in std_logic;
	green, yellow, red: out std_logic_vector(3 downto 0); output: integer);
end entity;

architecture Arch of TrafficLightContainer is
begin
			
	process(clk, rst)
	variable counter: integer range 0 to 6 := 0;
	variable current_lane: integer range 0 to 3 := 0;
	
	begin
		if rising_edge(clk) then
			output <= counter;
			if rst = '1' then
				counter :=  0;
				green <= "1000";
				yellow <= "0000";
				red <= "0111";
				current_lane := 0;
			end if;
			
			if counter = 5 then
--				green(current_lane) <= '0';
--				yellow(current_lane) <= '1';
				green <= "1000";
				yellow <= "0000";
				red <= "0111";
				counter := counter + 1;
				
			elsif counter = 6 then
--				yellow(current_lane) <= '0';
--				red(current_lane) <= '1';
				green <= "1000";
				yellow <= "0000";
				red <= "0111";
				
				
				if current_lane = 3 then
					current_lane := 0;
				else
					current_lane := current_lane + 1;
				end if;
--				red(current_lane) <= '0';
--				green(current_lane) <= '1';
				green <= "1000";
				yellow <= "0000";
				red <= "0111";
				counter := 0;
			else 
				counter := counter + 1;
			end if;
			
			
			
		end if;
	end process;
end Arch;
	