library ieee; 
use ieee.std_logic_1164.all;

entity OrFour is
	port ( x1,x2,x3,x4: std_logic;
	 R: out std_logic);
end entity;

architecture ARCH of OrFour is
	component OrGate is
		port (X,Y : in std_logic;
		O : out std_logic);
	end component;
	signal y1,y2: std_logic;
begin 
	Chip1: OrGate
		port map(x1, x2, y1);
	Chip2: OrGate
		port map(x3, x4, y2);
	Chip3: OrGate
		port map(y1, y2, R);
end;